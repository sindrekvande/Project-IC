*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../models/ptm_130_ngspice.spi
.include ../../lib/SUN_TR_GF130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6

VDD VDD VSS dc 1.5
VSS VSS 0 dc 0
VCOMP COMP VSS dc 0 PULSE(0, 1.5, 0, 10n, 10n, 30u, 60u, 0)
VIO IO VSS dc 0 PULSE(0, 1.5, 0, 10n, 10n, 29u, 60u, 0)
*VIO IO VSS dc 0 PULSE(0, 1.5, 0, 10n, 10n, 31u, 60u, 0) DATA low when comp. flips
VREAD READ VSS dc 0 PULSE(0, 1.5, 40u, 10n, 10n, 5u, 60u)

M4 DATA IO VDD VDD pmos w=0.5u  l=0.5u

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
.include cameraCircuit.cir
XDUT COMP DATA READ VSS MEMCELL

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set color0=white
set color1=black
unset askquit
tran 1n 60u

plot V(COMP) V(READ) V(DATA)

plot v(xdut.dmem) v(xdut.vg)
.endc
.end