
.SUBCKT PIXEL_SENSOR VBN1 VRAMP VRESET ERASE EXPOSE READ
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

XS1 VRESET VSTORE ERASE EXPOSE VDD VSS SENSOR

XC1 VCMP_OUT VSTORE VRAMP VBN1 VDD VSS COMP

XM1 READ VCMP_OUT DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS MEMORY

.ENDS
*///////////////////////////////////////////////////////////////////

.SUBCKT MEMORY READ VCMP_OUT
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

XM1 VCMP_OUT DATA_0 READ VSS MEMCELL
XM2 VCMP_OUT DATA_1 READ VSS MEMCELL
XM3 VCMP_OUT DATA_2 READ VSS MEMCELL
XM4 VCMP_OUT DATA_3 READ VSS MEMCELL
XM5 VCMP_OUT DATA_4 READ VSS MEMCELL
XM6 VCMP_OUT DATA_5 READ VSS MEMCELL
XM7 VCMP_OUT DATA_6 READ VSS MEMCELL
XM8 VCMP_OUT DATA_7 READ VSS MEMCELL

.ENDS
*///////////////////////////////////////////////////////////////////

.SUBCKT MEMCELL CMP DATA READ VSS
M12 VG CMP DATA VSS nmos  w=0.2u  l=0.13u
M13 DATA READ DMEM VSS nmos  w=0.4u  l=0.13u
M14 DMEM VG VSS VSS nmos  w=1u  l=0.13u
C2 VG VSS 1p
.ENDS
*///////////////////////////////////////////////////////////////////

.SUBCKT SENSOR VRESET VSTORE ERASE EXPOSE VDD VSS

C1 VSTORE VSS 100f
M1 VRESET ERASE VSTORE VSS nmos W=0.5u L=0.15u
M2 VPG EXPOSE VSTORE VSS nmos W=0.5u L=0.15u

Rphoto VPG VSS 1G
.ENDS
*///////////////////////////////////////////////////////////////////

.SUBCKT COMP VCMP_OUT VSTORE VRAMP VBN1 VDD VSS

M3 MGATE VSTORE BDRAIN VSS nmos W=0.5u L=0.15u
M4 BDRAIN VBN1 VSS VSS nmos W=0.5u L=0.15u
M5 MGATE MGATE VDD VDD pmos W={3.866*0.5u} L=0.15u
M6 RDRAIN MGATE VDD VDD pmos W={3.86*0.5u} L=0.15u
M7 RDRAIN VRAMP BDRAIN VSS nmos W=0.5u L=0.15u
M8 INODE RDRAIN VDD VDD pmos W={3.86*0.5u} L=0.15u
M9 INODE VBN1 VSS VSS nmos W=0.5u L=0.15u
M10 VCMP_OUT INODE VDD VDD pmos W={3.86*0.5u} L=0.15u
M11 VCMP_OUT INODE VSS VSS nmos W=0.5u L=0.15u

.ENDS
    