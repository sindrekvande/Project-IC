*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../models/ptm_130_ngspice.spi
.include ../../lib/SUN_TR_GF130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6

*----------------------------------------------------------------
* PARAMETERS
*----------------------------------------------------------------
.param TRF = 10n
.param TCLK = 100n
.param C_ERASE = 5
.param C_EXPOSE = 255
.param C_CONVERT = 255
.param C_READ = 5

*- Pulse Width of control signals
.param PW_ERASE =  {(C_ERASE +1)*TCLK}
.param PW_EXPOSE =  {(C_EXPOSE +1)*TCLK}
.param PW_CONVERT =  {(C_CONVERT +1)*TCLK}
.param PW_READ =  {(C_READ +1)*TCLK}

*- Delay of control signals
.param TD_ERASE = {TCLK }
.param TD_EXPOSE = {TD_ERASE + PW_ERASE + TCLK}
.param TD_CONVERT = {TD_EXPOSE + PW_EXPOSE + TCLK}
.param TD_READ = {TD_CONVERT + PW_CONVERT + TCLK}
.param PERIOD = {TD_READ + PW_READ + TCLK}

*- Analog parameters
.param VDD = 1.5
.param VADC_MIN = 0.5
.param VADC_MAX = 1.1
.param VADC_REF = {VADC_MAX - VADC_MIN}
.param VADC_LSB = {VADC_REF/256}

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
VDD VDD VSS dc VDD
VSS VSS 0 dc 0

*- Control signals
VERASE ERASE 0 dc 0 pulse (0 VDD TD_ERASE TRF TRF PW_ERASE PERIOD)
VEXPOSE EXPOSE 0 dc 0 pulse (0 VDD TD_EXPOSE TRF TRF PW_EXPOSE PERIOD)
VCONVERT CONVERT 0 dc 0 pulse (0 VDD TD_CONVERT TRF TRF PW_CONVERT PERIOD)
VREAD READ 0 dc 0 pulse (0 VDD TD_READ TRF TRF PW_READ PERIOD)

*- ADC related sources
VREF VREF 0 DC VADC_REF
VMAX VMAX 0 DC VADC_MAX
VRESET VRESET VMAX DC 0
VMIN VMIN 0 DC VADC_MIN

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
.include cameraCircuit.cir
XDUT READ VCMP_OUT 
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS MEMORY

VCMP_OUT VCMP_OUT VSS dc 0 PULSE(0, 1.5, 0, 10n, 10n, 35.8u, 53.4u, 0)

*----------------------------------------------------------------
* RAMP
*----------------------------------------------------------------
BR1 0 VRAMP I = V(CONVERT)*( 1n*(VADC_MAX - VADC_MIN)/PW_CONVERT)
CR1 VRAMP 0 1n ic=0

R1 VRAMP 0 1T

BR2 VRAMP VMIN I=V(ERASE)*V(VRAMP,VMIN)/100

*----------------------------------------------------------------
* Model the ramp generation and data for the memory
*----------------------------------------------------------------
B1 VADC 0 V = V(VRAMP) - VADC_MIN
XADC7 VADC   REST_7 VREF DATA_7  READ CONVERT VDD ADC_1BIT
XADC6 REST_7 REST_6 VREF DATA_6  READ CONVERT VDD ADC_1BIT
XADC5 REST_6 REST_5 VREF DATA_5  READ CONVERT VDD ADC_1BIT
XADC4 REST_5 REST_4 VREF DATA_4  READ CONVERT VDD ADC_1BIT
XADC3 REST_4 REST_3 VREF DATA_3  READ CONVERT VDD ADC_1BIT
XADC2 REST_3 REST_2 VREF DATA_2  READ CONVERT VDD ADC_1BIT
XADC1 REST_2 REST_1 VREF DATA_1  READ CONVERT VDD ADC_1BIT
XADC0 REST_1 REST_0 VREF DATA_0  READ CONVERT VDD ADC_1BIT
XDAC0 DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 DO VDD DAC_8BIT

*----------------------------------------------------------------
* 8-bit DAC model model
*----------------------------------------------------------------
* integer = 2^7*b7 + 2^6*b6 ... 2^0*b0
.SUBCKT DAC_8BIT DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 DO VDD
B1 DO_VDD 0 V=128*V(DATA_7)+64*V(DATA_6)+32*V(DATA_5)+16*V(DATA_4)+8*V(DATA_3)+4*V(DATA_2)+2*V(DATA_1)+1*V(DATA_0)
B2 DO 0 V = V(DO_VDD)/V(VDD)
.ENDS

*----------------------------------------------------------------
* 1-bit ADC model
*----------------------------------------------------------------
.SUBCKT ADC_1BIT VIN VOUT VREF DATA READ CONVERT VDD
B1 D 0 V= V(VIN) > V(VREF)/2 ? 1 : 0
B2 VOUT 0  V = 2*(V(VIN) - V(VREF)/2*V(D))
B3 DATA_INT 0 V = V(D)*V(VDD)
B4 DATA_INT DATA I=V(CONVERT)*V(DATA_INT,DATA)/1k
B5 DATA VDD I=V(READ)*V(DATA,VDD)/1e4
.ENDS

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set color0=white
set color1=black
unset askquit
tran 1n 60u

*plot V(DATA_0) V(XDUT.XM1.DMEM) V(VCMP_OUT) V(READ)
*plot V(DATA_1) V(XDUT.XM2.DMEM) V(VCMP_OUT) V(READ)
*plot V(DATA_2) V(XDUT.XM3.DMEM) V(VCMP_OUT) V(READ)
*plot V(DATA_3) V(XDUT.XM4.DMEM) V(VCMP_OUT) V(READ)
plot V(DATA_4) V(XDUT.XM5.DMEM) V(VCMP_OUT) V(READ)
plot V(DATA_5) V(XDUT.XM6.DMEM) V(VCMP_OUT) V(READ)
plot V(DATA_6) V(XDUT.XM7.DMEM) V(VCMP_OUT) V(READ)
plot V(DATA_7) V(XDUT.XM8.DMEM) V(VCMP_OUT) V(READ)

*plot V(XDUT.XM1.VG) V(XDUT.XM1.DMEM) V(VCMP_OUT) V(READ)
*plot V(XDUT.XM2.VG) V(XDUT.XM2.DMEM) V(VCMP_OUT) V(READ) 
*plot V(XDUT.XM3.VG) V(XDUT.XM3.DMEM) V(VCMP_OUT) V(READ)
*plot V(XDUT.XM4.VG) V(XDUT.XM4.DMEM) V(VCMP_OUT) V(READ) 
*plot V(XDUT.XM5.VG) V(XDUT.XM5.DMEM) V(VCMP_OUT) V(READ)
*plot V(XDUT.XM6.VG) V(XDUT.XM6.DMEM) V(VCMP_OUT) V(READ) 
*plot V(XDUT.XM7.VG) V(XDUT.XM7.DMEM) V(VCMP_OUT) V(READ)
*plot V(XDUT.XM8.VG) V(XDUT.XM8.DMEM) V(VCMP_OUT) V(READ) 
.endc
.end