*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../models/ptm_130_ngspice.spi
.include ../../lib/SUN_TR_GF130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6


*evt. bruke pmos inn til data???
*-> Sikkert ikke nødvendig for våres del, men fint å ha hvis man ønsker å brife litt?

*----------------------------------------------------------------
* PARAMETERS
*----------------------------------------------------------------

.param TRF = 10n
.param TCLK = 100n
.param C_ERASE = 5
.param C_EXPOSE = 255
.param C_CONVERT = 255
.param C_READ = 5

*- Pulse Width of control signals
.param PW_ERASE =  {(C_ERASE +1)*TCLK}
.param PW_EXPOSE =  {(C_EXPOSE +1)*TCLK}
.param PW_CONVERT =  {(C_CONVERT +1)*TCLK}
.param PW_READ =  {(C_READ +1)*TCLK}

*- Delay of control signals
.param TD_ERASE = {TCLK }
.param TD_EXPOSE = {TD_ERASE + PW_ERASE + TCLK}
.param TD_CONVERT = {TD_EXPOSE + PW_EXPOSE + TCLK}
.param TD_READ = {TD_CONVERT + PW_CONVERT + TCLK}
.param PERIOD = {TD_READ + PW_READ + TCLK}

*- Analog parameters
.param VDD = 1.5
.param VADC_MIN = 0.5
.param VADC_MAX = 1.1
.param VADC_REF = {VADC_MAX - VADC_MIN}
.param VADC_LSB = {VADC_REF/256}

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
VDD VDD VSS dc VDD
VSS VSS 0 dc 0

*- Control signals
VREAD READ 0 dc 0 pulse (0 VDD TD_READ TRF TRF PW_READ PERIOD)
VCONVERT CONVERT 0 dc 0 pulse (0 VDD TD_CONVERT TRF TRF PW_CONVERT PERIOD)

*- ADC related sources
VREF VREF 0 DC VADC_REF
VMAX VMAX 0 DC VADC_MAX
*VRESET VRESET VMAX DC 0
VMIN VMIN 0 DC VADC_MIN

**----------------------------------------------------------------
** DUT
*----------------------------------------------------------------
.include cameraCircuit.cir
XDUT VRESET VSTORE ERASE EXPOSE VDD VSS SENSOR
XDUT VCMP_OUT VSTORE VRAMP VBN1 VDD VSS COMP
XDUT COMP DATA READ VSS MEMCELL

*----------------------------------------------------------------
* 1-bit ADC model
*----------------------------------------------------------------
* Model the DATA output as pulled to VDD when we're reading
.SUBCKT ADC_1BIT VIN VOUT VREF DATA READ CONVERT VDD
B1 D 0 V= V(VIN) > V(VREF)/2 ? 1 : 0
B2 VOUT 0  V = 2*(V(VIN) - V(VREF)/2*V(D))
B3 DATA_INT 0 V = V(D)*V(VDD)
B4 DATA_INT DATA I=V(CONVERT)*V(DATA_INT,DATA)/1k
B5 DATA VDD I=V(READ)*V(DATA,VDD)/1e4
.ENDS


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------

.control
set color0=white
set color1=black
unset askquit
tran 1n 60u

plot V(COMP) V(READ) V(DATA)

plot v(xdut.xm1.xm1.vg) v(xdut.xm1.xm1.dmem)
plot v(xdut.xm1.xm2.vg) v(xdut.xm1.xm2.dmem)
plot v(xdut.xm1.xm3.vg) v(xdut.xm1.xm3.dmem)
plot v(xdut.xm1.xm4.vg) v(xdut.xm1.xm4.dmem)
plot v(xdut.xm1.xm5.vg) v(xdut.xm1.xm5.dmem)
plot v(xdut.xm1.xm6.vg) v(xdut.xm1.xm6.dmem)
plot v(xdut.xm1.xm7.vg) v(xdut.xm1.xm7.dmem)
plot v(xdut.xm1.xm8.vg) v(xdut.xm1.xm8.dmem)
.endc
.end